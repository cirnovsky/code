module sl
